library verilog;
use verilog.vl_types.all;
entity counter_bonus_tb is
end counter_bonus_tb;
