library verilog;
use verilog.vl_types.all;
entity counter8bit_tb is
end counter8bit_tb;
